// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
    parameter BITS = 32
) (
`ifdef USE_POWER_PINS
    inout vdda1,	// User area 1 3.3V supply
    inout vdda2,	// User area 2 3.3V supply
    inout vssa1,	// User area 1 analog ground
    inout vssa2,	// User area 2 analog ground
    inout vccd1,	// User area 1 1.8V supply
    inout vccd2,	// User area 2 1.8v supply
    inout vssd1,	// User area 1 digital ground
    inout vssd2,	// User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
    inout [`MPRJ_IO_PADS-10:0] analog_io,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

/*--------------------------------------*/
/* User project is instantiated  here   */
/*--------------------------------------*/


SRAM_Wrapper_top SRAM_IMC_TOP(

.clk(wb_clk_i),					//Common clock
.reset_n(wb_rst_i),					//wb_rst_i	
.wbs_we_i(wbs_we_i) ,					//wbs_we_i=0 for read ;wbs_we_i=1 for write		
.wishbone_buffer_data_in(wbs_dat_i), 			//wbs_dat_i
.wishbone_rw_addr(wbs_adr_i),				//wishbone_addr
.wishbone_databus_out(wbs_dat_o),	 		//wbs_dat_o
.VCLP(analog_io[11]),					// connect to Analog IO
.EN(analog_io[12]),					// connect to Analog IO
.Iref0(analog_io[7]),					// connect to Analog IO
.Iref1(analog_io[8]),					// connect to Analog IO
.Iref2(analog_io[9]),					// connect to Analog IO
.Iref3(analog_io[13]),					// connect to Analog IO
.Iout0(analog_io[14]),					// Deepak -30/12/22 - added for MPW8
.Iout1(analog_io[15]),					// Deepak -30/12/22 - added for MPW8
.Iout2(analog_io[16]),					// Deepak -30/12/22 - added for MPW8
.Iout3(analog_io[17]),					// Deepak -30/12/22 - added for MPW8
.EN_VCLP(la_data_out[0]),				//Deepak_28/11/22: needs to be passed to analog DUT for EN & VCLP enable
.MAC_starting(la_data_out[1]),				// Deepak : Enable for MUX for Iref			
.OB_demux(la_data_out[2]),				// Deepak: select line for Irefs
.controller_opcode(la_data_out[5:3]),
.controller_ext_state(la_data_out[7:6]),
.controller_int_state(la_data_out[10:8]),
.full_IB(la_data_out[11]),
.full_WB(la_data_out[12]), 
.full_SA(la_data_out[13]), 
.full_OB(la_data_out[14]),
.empty_IB(la_data_out[15]), 
.empty_WB(la_data_out[16]), 
.empty_SA(la_data_out[17]), 
.empty_OB(la_data_out[18])
); 




/*

user_proj_example mprj (
`ifdef USE_POWER_PINS
	.vccd1(vccd1),	// User area 1 1.8V power
	.vssd1(vssd1),	// User area 1 digital ground
`endif

    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),

    // MGMT SoC Wishbone Slave

    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .wbs_sel_i(wbs_sel_i),
    .wbs_adr_i(wbs_adr_i),
    .wbs_dat_i(wbs_dat_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_dat_o(wbs_dat_o),

    // Logic Analyzer

    .la_data_in(la_data_in),
    .la_data_out(la_data_out),
    .la_oenb (la_oenb),

    // IO Pads

    .io_in (io_in),
    .io_out(io_out),
    .io_oeb(io_oeb),

    // IRQ
    .irq(user_irq)
);

*/

endmodule	// user_project_wrapper

`default_nettype wire
